��   ��A��*SYST�EM*��V7.7�079 3/2�7/2013 �A   ����AW_SCH_�T   � �$CMD_VOLkTS 6WF?�AMP?PKU
F�REQYULSE�@SPEED@T{IM�FDBK:��UOMMENT� & SA�DVISE- ` �%6�;�U
I	bt�$�$CLASS  ����J��~���$AWE* � R J��  @ �<A�  B� �w��@�BH��N�NCo�)Q��|a�p������?�����	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o�o�o�o +=Oas��� ������'�9� K�]�o���������ɋ���Runinx����=���߆�	 Burnba�ck.�@�R�  Wirestih��S�@،Ӂ��� OnTheFly� �u�"�p���S�e�+� =�������ǟٟ럍 ��c��C�U��-� �������ɯۯ�� �P�ں3�E���{� ��۵����˿�D�� @���#�5����k�}� �ŗϩϻϽ�5��� 1߻��%�����[�m� �Շߙ߽߫�%��� !��������K�]� ��w��������� ���������;�M���pg�y�[� 2fo @%��tti �: T=0.8 �W�S=10 C�O2=15�B���}،�
1.0D���}��2�I9���6� �'1� L�2D�m55�Ћ�4���3(�20|�r��f��4.5����"\-Filglet�4C��A�Z*�y+���/ �()�K�/�.i�$�1��Z*�9;��#CRL?^&�24�����?^&')�=�v� C�-Lapi b*�/ B��OG�/�C!�!�LO^H)8ptOׁJH2.3�O
<(����O�Lm�I � _��CA�H?J�'/yK�1z-C-J�oint�Ou_�� �_�V�O�[�A�Xg_ ���RK^�X�_�0F?  